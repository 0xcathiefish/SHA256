`timescale  1ns/1ns

module sha256_tb;

    parameter cycle = 2;

    reg clk,rst;

    reg [511:0] cin;

    //reg [3:0]   cmd_state;

    wire [255:0] out;




Sha256 Sha_1(clk,rst,cin,out);

initial begin

    rst = 1;
    clk = 1;

    forever begin
        
        #(cycle/2) clk = ~clk;
    end
end

initial begin

    cin = 0;
    //cmd_state = 0;
end


initial begin

    #10;

    rst <= 0;

    cin <= 512'h696C6F76657580000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030;


    //cmd_state = 4'd1;


end


endmodule


// 01101001011011000110111101110110011001010111010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000